////////////////////////////////////////////////////////////////////////////////
// @file    tb_converter.v
// @author  JAY CONVERTINO
// @date    2021.06.21
// @brief   UTIL AXIS DATA WIDTH CONVERTER
////////////////////////////////////////////////////////////////////////////////

`timescale 1 ns/10 ps

module tb_converter;
  
  reg         tb_data_clk = 0;
  reg         tb_rst = 0;
  //master
  wire [15:0] tb_dmaster;
  wire        tb_vmaster;
  reg         tb_rmaster;
  //slave
  reg [127:0] tb_dslave;
  reg         tb_vslave;
  wire        tb_rslave;
  reg         tb_vslave_off;
  reg         tb_vslave_toggle = 0;
  
  
  
  localparam CLK_PERIOD = 500;
  localparam RST_PERIOD = 1000;
  
  util_axis_data_width_converter #(
    .master_width(2),
    .slave_width(16)
  ) dut (
    //axi streaming clock and reset.
    .aclk(tb_data_clk),
    .arstn(~tb_rst),
    //1553
    //master data out interface
    .m_axis_tdata(tb_dmaster),
    .m_axis_tvalid(tb_vmaster),
    .m_axis_tready(tb_rmaster),
    //slave data in interface
    .s_axis_tdata(tb_dslave),
    .s_axis_tvalid(tb_vslave),
    .s_axis_tready(tb_rslave)
  );
    
  //reset
  initial
  begin
    tb_rst <= 1'b1;
    tb_vslave_off <= 1'b1;
    
    #RST_PERIOD;
    
    tb_rst <= 1'b0;
    
    #30000;
    
    tb_vslave_off <= 1'b0;
    
    #30500;
    
    tb_vslave_off <= 1'b1;
  end
  
  //copy pasta, vcd generation
  initial
  begin
    $dumpfile("sim/icarus/tb_converter.vcd");
    $dumpvars(0,tb_converter);
  end
  
  //clock
  always
  begin
    tb_data_clk <= ~tb_data_clk;
    
    #(CLK_PERIOD/4);
  end
  
  //valid off/on
  always
  begin
    tb_vslave_toggle <= ~tb_vslave_toggle;
    
    #(CLK_PERIOD/2);
  end
  
  //product data
  always @(posedge tb_data_clk)
  begin
    if (tb_rst == 1'b1) begin
      tb_dslave <= 128'h55005500550055005500550055005500;
      tb_vslave <= 0;
      tb_rmaster<= 0;
    end else begin
      tb_rmaster  <= $random % 2;
      tb_vslave   <= tb_vslave_off;
      
      tb_dslave   <= tb_dslave;
      
      if((tb_rslave == 1'b1) && (tb_vslave_off == 1'b1)) begin
        tb_dslave <= tb_dslave + 128'h01010101010101010101010101010101;
      end
    end
  end
  
  //copy pasta, no way to set runtime... this works in vivado as well.
  initial begin
    #1_000_000; // Wait a long time in simulation units (adjust as needed).
    $display("END SIMULATION");
    $finish;
  end
endmodule

